module STORED_IMAGES_DECODER (CLM, ROW, IMG_ID, COLOR);

	input logic  [4:0] CLM, ROW;
	input logic  [9:0] IMG_ID;
	output logic [3:0] COLOR;
	logic [3:0] SPRITE [0:31][0:31];
	assign SPRITE =
	'{'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0011, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0011, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0001, 4'b0000, 4'b0011, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0011, 4'b0001, 4'b0000, 4'b0001, 4'b0000, 4'b0011, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0001, 4'b0000, 4'b0001, 4'b0001, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0011, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0000, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0000, 4'b0001, 4'b0000, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b0011, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0100, 4'b0100, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0100, 4'b0100, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},'{  
		4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}
	};
	
	assign COLOR = SPRITE [CLM][ROW];

endmodule 