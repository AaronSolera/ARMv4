module NEW_INSTRUCTION_VERIFICATOR (HF_CLK, RST, INSTRUCTION, NOT_EQU);
	
	input logic HF_CLK, RST;
	input logic [31:0] INSTRUCTION;
	output logic NOT_EQU;
	logic W_EQU;
	logic [31:0] OLD_INSTRUCTION;
	
	EQUAL_COMPARATOR_MODULE #(32) 
		EQU_CMP (INSTRUCTION, OLD_INSTRUCTION, W_EQU);
		
	REGISTER_MODULE #(32)
		MM (HF_CLK, RST, ~W_EQU, INSTRUCTION, OLD_INSTRUCTION);

	assign NOT_EQU = ~W_EQU;
		 
endmodule 