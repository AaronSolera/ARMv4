module GRAPHIC_PROCESSING_UNIT (CLK, RST, INSTRUCTION, H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, R, G, B);
	
	input  logic CLK, RST;
	input  logic [31:0] INSTRUCTION;
	output logic H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N;
	output logic [7:0] R, G, B;
	
	logic ENA_BACKGROUND_COLOR;
	logic [9:0]  SCREEN_POS_X, SCREEN_POS_Y;
	logic [15:0] CURRENT_INSTRUCTION;
	logic [3:0]  ID_COLOR, IMG_COLOR;
	logic [23:0] RGB_COLOR;
	
	VGA_CONTROLLER_MODULE 
		VGA_CM (CLK, RST, H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, SCREEN_POS_X, SCREEN_POS_Y);
	 
	GRAPHIC_INSTRUCTION_CONTROL_UNIT 
		GICU (CLK, RST, SCREEN_POS_X, SCREEN_POS_Y, {10'd0, 10'd0, 12'd0}, CURRENT_INSTRUCTION);
		
	STORED_IMAGES_DECODER 
		SID (CURRENT_INSTRUCTION[4:0], CURRENT_INSTRUCTION[9:5], CURRENT_INSTRUCTION[15:10], IMG_COLOR);
	
	N_INPUTS_AND #(6)
		BACKGROUND_COLOR (CURRENT_INSTRUCTION[15:10],ENA_BACKGROUND_COLOR);
		
	N_BITS_ONE_SELECT_MUX_MODULE #(4)
		COLOR_MUX (IMG_COLOR, 4'hF, ENA_BACKGROUND_COLOR, ID_COLOR);

	COLOR_DECODER 
		CD (ID_COLOR, RGB_COLOR);
	
	assign R = RGB_COLOR[23:16];
	assign G = RGB_COLOR[15:8];
	assign B = RGB_COLOR[7:0];
	
endmodule 