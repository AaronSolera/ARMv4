module DECODER_UNIT(input logic [5:0] Funct, input logic [1:0] Op, input logic [3:0] Rd);
	//Main Decoder
	//PC Logic
	//ALU Logic
endmodule