module STORED_IMAGES_DECODER (CLM, ROW, IMG_ID, COLOR);

	input logic  [4:0] CLM, ROW;
	input logic  [9:0] IMG_ID;
	output logic [3:0] COLOR;
	logic [3:0] SPRITE [0:1][0:31][0:31];
	assign SPRITE =
	'{
		'{
		'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b000, 3'b001, 3'b001, 3'b010},'{ 
		3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b010, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b011, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b011, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b011, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b011, 3'b001, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b011, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001
		}
		},
		'{
		'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b000, 3'b001, 3'b001, 3'b010},'{ 
		3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b010, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b011, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b011, 3'b011, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b011, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b011, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b010, 3'b001, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b010, 3'b010, 3'b011, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b011, 3'b001, 3'b000, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b000, 3'b011, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001},'{ 
		3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001
		}
		}
	};
	assign COLOR = SPRITE [IMG_ID][CLM][ROW];

endmodule 