module GRAPHIC_CONTROL_UNIT (HF_CLK, RST, INS, BLANK, CURRENT_INS, SID_CLM, SID_ROW, PGA_CLM, PGA_ROW);

	input  logic        HF_CLK, RST, BLANK;
	input  logic [31:0] INS;
	output logic [9:0]  PGA_CLM, PGA_ROW;
	output logic [4:0]  SID_CLM, SID_ROW;
	output logic [31:0] CURRENT_INS;
	
	logic SID_CLM_CLK, SID_ROW_CLK, PGA_CLM_COUT, PGA_ROW_COUT, INVISIBLE_INS, INS_CMLPTED, CHANGE_C_INS;
	logic [4:0] W_SID_CLM, W_SID_ROW;
	logic [31:0] C_INS;
	
	INSTRUCTION_CONTROL_UNIT 
		ICU (HF_CLK, RST, BLANK, CHANGE_C_INS, INS, C_INS);
	
	COUNTER_MODULE 
		SID_CLM_CM  (HF_CLK,      BLANK & RST, W_SID_CLM),
		SID_ROW_CM  (SID_CLM_CLK, BLANK & RST, W_SID_ROW);
		
	EQUAL_COMPARATOR_MODULE #(5)
		SID_CLM_CMP (W_SID_CLM, 5'd32, SID_CLM_CLK),
		SID_ROW_CMP (W_SID_ROW, 5'd32, SID_ROW_CLK);
	EQUAL_COMPARATOR_MODULE #(3)
		INVISIBLE_INS_CMP (C_INS[12:10], 3'b111, INVISIBLE_INS);
	
	ADDER_MODULE #(10) 
		PGA_CLM_ADDER (W_SID_CLM, C_INS[31:22], 1'b0, PGA_CLM, PGA_CLM_COUT),
		PGA_ROW_ADDER (W_SID_ROW, C_INS[21:13], 1'b0, PGA_ROW, PGA_ROW_COUT);
	
	_AND
		AND (SID_CLM_CLK, SID_ROW_CLK, INS_CMLPTED);
		
	_OR
		INVISIBLE_OR (INS_CMLPTED, INVISIBLE_INS, CHANGE_C_INS);
	
	assign SID_CLM = W_SID_CLM;
	assign SID_ROW = W_SID_ROW;
	assign CURRENT_INS = C_INS;
	
endmodule 