module NEW_INSTRUCTION_VERIFICATOR (HF_CLK, RST, INSTRUCTION, EQU, NOT_EQU);
	
	input logic HF_CLK, RST;
	input logic [31:0] INSTRUCTION;
	output logic EQU, NOT_EQU;
	logic W_EQU;
	logic [31:0] OLD_INSTRUCTION;
	
	REGISTER_MODULE #(32)
		MM (HF_CLK, RST, ~W_EQU, INSTRUCTION, OLD_INSTRUCTION);
	
	EQUAL_COMPARATOR_MODULE #(32) 
		EQU_CMP (INSTRUCTION, OLD_INSTRUCTION, W_EQU);
		
	assign EQU = W_EQU;
	assign NOT_EQU = ~W_EQU;
		
endmodule 