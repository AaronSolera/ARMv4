module GRAPHIC_INSTRUCTION_CONTROL_UNIT (CLK, RST, SYS_X, SYS_Y, INS, C_INS);

	input  logic        CLK, RST;
	input  logic [9:0]  SYS_X, SYS_Y;
	input  logic [31:0] INS;
	output logic [15:0] C_INS;
	logic WRITE;
	
	logic [5:0] NEW_INS_ADD;
	logic CYCLE_X_RST, CYCLE_Y_RST, SYS_RST, MASTER_RST;

	EQUAL_COMPARATOR_MODULE #(10)
		SYS_X_RESET (SYS_X, 10'd634, CYCLE_X_RST),
		SYS_Y_RESET (SYS_Y, 10'd479, CYCLE_Y_RST);

	_AND
		SYS_RST_AND (CYCLE_X_RST, CYCLE_Y_RST, SYS_RST),
		MASTER_RST_AND (~SYS_RST, RST, MASTER_RST);
		
	NEW_INSTRUCTION_VERIFICATOR 
		NIV (CLK, MASTER_RST, INS, WRITE);      
	
	COUNTER_MODULE 
		NEW_INS_CM  (~WRITE, MASTER_RST, NEW_INS_ADD);
	
	GRAPHIC_INSTRUCTION_MEMORY_MODULE
		GRAPHIC_INSTRUCTION_MEMORY (CLK, MASTER_RST, SYS_X, SYS_Y, NEW_INS_ADD, WRITE, INS, C_INS);
		
endmodule 