module EIGHT_N_BITS_INPUTS_THREE_BITS_SELECT_MUX_MODULE #(parameter BITS = 3) (DATA, SELECT, OUT);

	input logic [7:0][BITS-1:0] DATA;
	input logic [2:0] SELECT;
	output logic [BITS-1:0] OUT;
	logic [BITS-1:0] W_FIRST_MUX, W_SECOND_MUX;
	
	FOUR_N_BITS_INPUTS_TWO_BITS_SELECT_MUX_MODULE #(BITS)
		FIRST_MUX (DATA[3:0], SELECT[1:0], W_FIRST_MUX),
		SECOND_MUX (DATA[7:4], SELECT[1:0], W_SECOND_MUX);
	N_BITS_ONE_SELECT_MUX_MODULE #(BITS)
		THIRD_MUX (W_FIRST_MUX, W_SECOND_MUX, SELECT[2], OUT);
	
endmodule 