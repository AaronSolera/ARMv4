module AREA_VERIFICATOR_MODULE (X, Y, POS_X, POS_Y, DIFF_X_COUNT, DIFF_Y_COUNT, IN_AREA_INDICATOR);

	input logic [9:0] POS_X, X, POS_Y, Y;
	output logic IN_AREA_INDICATOR;
	output logic [4:0] DIFF_X_COUNT, DIFF_Y_COUNT;
	logic [9:0] POSX_MIN_X, POSY_MIN_Y, POSX_MIN_XW, POSY_MIN_YH;
	logic GTX, LTXW, GTY, LTYH, X_AREA_INDICATOR, Y_AREA_INDICATOR;
		
	FULL_N_BITS_SUBTRACTOR_MODULE #(10) 
		POSX_GT_X  (POS_X, X, POSX_MIN_X, GTX),
		POSY_GT_Y  (POS_Y, Y, POSY_MIN_Y, GTY),
		POSX_LT_XW (10'd31, POSX_MIN_X, POSX_MIN_XW, LTXW),
		POSY_LT_YH (10'd31, POSY_MIN_Y, POSY_MIN_YH, LTYH);
		
	_NOR
		X_AREA_NOR (GTX, LTXW, X_AREA_INDICATOR),
		Y_AREA_NOR (GTY, LTYH, Y_AREA_INDICATOR);
		
	_AND AND (X_AREA_INDICATOR, Y_AREA_INDICATOR, IN_AREA_INDICATOR); 
	
	assign DIFF_X_COUNT = POSX_MIN_X[4:0];
	assign DIFF_Y_COUNT = POSY_MIN_Y[4:0];
	
endmodule  