module SIXTEEN_N_BITS_INPUTS_FOUR_BITS_SELECT_MUX_MODULE #(parameter BITS = 3) (DATA, SELECT, OUT);

	input logic [15:0][BITS-1:0] DATA;
	input logic [3:0] SELECT;
	output logic [BITS-1:0] OUT;
	logic [BITS-1:0] W_FIRST_MUX, W_SECOND_MUX;
	
	EIGHT_N_BITS_INPUTS_THREE_BITS_SELECT_MUX_MODULE #(BITS)
		FIRST_MUX (DATA[7:0], SELECT[2:0], W_FIRST_MUX),
		SECOND_MUX (DATA[15:8], SELECT[2:0], W_SECOND_MUX);
	N_BITS_ONE_SELECT_MUX_MODULE #(BITS)
		THIRD_MUX (W_FIRST_MUX, W_SECOND_MUX, SELECT[3], OUT);
	
endmodule 