module GRAPHIC_PROCESSING_UNIT (CLK, RST, INSTRUCTION, H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, RGB_COLOR);
	
	//Instruction = Y[10],X[10],OP[3],SPRITE_ID[9]
	input  logic        CLK, RST;
	input  logic [31:0] INSTRUCTION;
	output logic        H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N;
	output logic [23:0] RGB_COLOR; 
	
	logic        REFRESH;
	logic [31:0] CURRENT_INSTRUCTION;
	logic [9:0]  PGA_CLM, PGA_ROW, SCREEN_POS_X, SCREEN_POS_Y, PGA_CLM_MUX, PGA_ROW_MUX;
	logic [4:0]  SID_CLM, SID_ROW;
	logic [3:0]  SID_COLOR;
	
	VGA_CONTROLLER_MODULE 
		VCM (CLK, RST, H_SYNC, REFRESH, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, SCREEN_POS_X, SCREEN_POS_Y);
	
	GRAPHIC_CONTROL_UNIT 
		GCU (CLK, RST, INSTRUCTION, REFRESH, CURRENT_INSTRUCTION, SID_CLM, SID_ROW, PGA_CLM, PGA_ROW);

	N_BITS_ONE_SELECT_MUX_MODULE #(10)
		PGA_CLM_MUX_MODULE (PGA_CLM, SCREEN_POS_X, REFRESH, PGA_CLM_MUX),
		PGA_ROW_MUX_MODULE (PGA_ROW, SCREEN_POS_Y, REFRESH, PGA_ROW_MUX);
	
	STORED_IMAGES_DECODER SID (SID_CLM, SID_ROW, CURRENT_INSTRUCTION[9:0], SID_COLOR);
	
	PIXEL_GRAPHIC_ARRAY #(4) 
		PGA (CLK, RST, ~REFRESH, PGA_ROW_MUX, PGA_CLM_MUX, SID_COLOR, RGB_COLOR);
	
	assign V_SYNC = REFRESH;
	
endmodule 