module VGA_CONTROLLER_MODULE (CLK, RST, H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, SCREEN_POS_X, SCREEN_POS_Y);
	
	input logic CLK, RST;
	output logic H_SYNC, V_SYNC, VGA_CLK, VGA_SYNC_N, VGA_BLANK_N;
	output logic [9:0] SCREEN_POS_X, SCREEN_POS_Y;
	logic OUT_CLK, H_CLK, V_CLK, H_RGB_ENA, V_RGB_ENA;
	
	CLK_HALF_DIV_MODULE 
		F_DIV (CLK, RST, OUT_CLK);
		
	SYNC_MODULE 
		H_SYNC_MODULE (OUT_CLK, RST, 10'd95, 10'd143, 10'd778, 10'd793, H_RGB_ENA, H_CLK, SCREEN_POS_X),
		V_SYNC_MODULE (H_CLK,   RST, 10'd2,  10'd35,  10'd515, 10'd524, V_RGB_ENA, V_CLK, SCREEN_POS_Y);
	
	_AND
		VGA_SYNC_AND  (H_CLK,     V_CLK,     VGA_SYNC_N),
		VGA_BLANK_AND (H_RGB_ENA, V_RGB_ENA, VGA_BLANK_N);
		
	assign H_SYNC  =  H_CLK;
	assign V_SYNC  =  V_CLK;
	assign VGA_CLK =  OUT_CLK;
	
endmodule 