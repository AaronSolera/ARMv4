module INSTRUCTION_CONTROL_UNIT (HF_CLK, RST, BLANK, CHANGE_C_INS, INS, C_INS);

	input  logic        HF_CLK, BLANK, RST, CHANGE_C_INS;
	input  logic [31:0] INS;
	output logic [31:0] C_INS;
	logic WRITE;
	
	logic [9:0] NEW_INS_ADD, READ_INS_ADD, GIM_ADD;
	logic ALL_INS_CMLPTED, EQU;
	
	NEW_INSTRUCTION_VERIFICATOR 
		NIV (HF_CLK, ~BLANK & RST, INS, EQU, WRITE);
		
	COUNTER_MODULE 
		NEW_INS_CM  (WRITE,        ~BLANK & RST, NEW_INS_ADD),
		READ_INS_CM (CHANGE_C_INS, ~BLANK & RST, READ_INS_ADD);
		
	N_BITS_ONE_SELECT_MUX_MODULE #(10)
		INS_ADD_MUX (READ_INS_ADD, NEW_INS_ADD, WRITE, GIM_ADD);
	
	MEMORY_MODULE #(32, 10)
		GRAPHIC_INSTRUCTION_MEMORY (~HF_CLK, ~BLANK & RST, GIM_ADD, WRITE, INS, C_INS);
		
endmodule 